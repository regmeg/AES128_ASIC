`line 1 "verilog/v_hier_noport.v" 0
// DESCRIPTION: Verilog-Perl: Example Verilog for testing package
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2000-2012 by Wilson Snyder.

module v_hier_noport;
   reg internal;
endmodule
