`line 1 "verilog/t_86_vhier_tick_sub.v" 0
// DESCRIPTION: Verilog::Preproc: Example source code
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2000-2012 by Wilson Snyder.

module t_86_vhier_tick_sub;
endmodule
